module rr_arb (
              input clk,
              input rst_n,
              input [2:0] req,
              output logic [2:0]  grant
);
 
